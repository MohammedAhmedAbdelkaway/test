

// First.
module wire
{
input x,
output y};

assign y = x;

endmodule